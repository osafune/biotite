// nios2core.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module nios2core (
		input  wire        clk_clk,         //     clk.clk
		inout  wire [11:0] gpio0_export,    //   gpio0.export
		inout  wire [11:0] gpio1_export,    //   gpio1.export
		inout  wire [11:0] gpio2_export,    //   gpio2.export
		output wire [23:0] led7seg_export,  // led7seg.export
		inout  wire [3:0]  qspi_sio,        //    qspi.sio
		output wire        qspi_sck,        //        .sck
		output wire        qspi_ce_n,       //        .ce_n
		input  wire        qspi_outclock,   //        .outclock
		input  wire        reset_reset_n,   //   reset.reset_n
		input  wire [2:0]  syskey_in_port,  //  syskey.in_port
		output wire [2:0]  syskey_out_port  //        .out_port
	);

	wire  [31:0] nios2_e_data_master_readdata;                                        // mm_interconnect_0:nios2_e_data_master_readdata -> nios2_e:d_readdata
	wire         nios2_e_data_master_waitrequest;                                     // mm_interconnect_0:nios2_e_data_master_waitrequest -> nios2_e:d_waitrequest
	wire         nios2_e_data_master_debugaccess;                                     // nios2_e:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_e_data_master_debugaccess
	wire  [28:0] nios2_e_data_master_address;                                         // nios2_e:d_address -> mm_interconnect_0:nios2_e_data_master_address
	wire   [3:0] nios2_e_data_master_byteenable;                                      // nios2_e:d_byteenable -> mm_interconnect_0:nios2_e_data_master_byteenable
	wire         nios2_e_data_master_read;                                            // nios2_e:d_read -> mm_interconnect_0:nios2_e_data_master_read
	wire         nios2_e_data_master_write;                                           // nios2_e:d_write -> mm_interconnect_0:nios2_e_data_master_write
	wire  [31:0] nios2_e_data_master_writedata;                                       // nios2_e:d_writedata -> mm_interconnect_0:nios2_e_data_master_writedata
	wire  [31:0] nios2_e_instruction_master_readdata;                                 // mm_interconnect_0:nios2_e_instruction_master_readdata -> nios2_e:i_readdata
	wire         nios2_e_instruction_master_waitrequest;                              // mm_interconnect_0:nios2_e_instruction_master_waitrequest -> nios2_e:i_waitrequest
	wire  [27:0] nios2_e_instruction_master_address;                                  // nios2_e:i_address -> mm_interconnect_0:nios2_e_instruction_master_address
	wire         nios2_e_instruction_master_read;                                     // nios2_e:i_read -> mm_interconnect_0:nios2_e_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;              // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;           // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_readdata;      // peridot_qspi_psram_0:avs_readdata -> mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_waitrequest;   // peridot_qspi_psram_0:avs_waitrequest -> mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_waitrequest
	wire  [22:0] mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_address;       // mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_address -> peridot_qspi_psram_0:avs_address
	wire         mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_read;          // mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_read -> peridot_qspi_psram_0:avs_read
	wire   [3:0] mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_byteenable;    // mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_byteenable -> peridot_qspi_psram_0:avs_byteenable
	wire         mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_readdatavalid; // peridot_qspi_psram_0:avs_readdatavalid -> mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_write;         // mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_write -> peridot_qspi_psram_0:avs_write
	wire  [31:0] mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_writedata;     // mm_interconnect_0:peridot_qspi_psram_0_avalon_slave_0_writedata -> peridot_qspi_psram_0:avs_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                      // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                       // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_boot_flash_csr_readdata;                           // boot_flash:avmm_csr_readdata -> mm_interconnect_0:boot_flash_csr_readdata
	wire   [0:0] mm_interconnect_0_boot_flash_csr_address;                            // mm_interconnect_0:boot_flash_csr_address -> boot_flash:avmm_csr_addr
	wire         mm_interconnect_0_boot_flash_csr_read;                               // mm_interconnect_0:boot_flash_csr_read -> boot_flash:avmm_csr_read
	wire         mm_interconnect_0_boot_flash_csr_write;                              // mm_interconnect_0:boot_flash_csr_write -> boot_flash:avmm_csr_write
	wire  [31:0] mm_interconnect_0_boot_flash_csr_writedata;                          // mm_interconnect_0:boot_flash_csr_writedata -> boot_flash:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_boot_flash_data_readdata;                          // boot_flash:avmm_data_readdata -> mm_interconnect_0:boot_flash_data_readdata
	wire         mm_interconnect_0_boot_flash_data_waitrequest;                       // boot_flash:avmm_data_waitrequest -> mm_interconnect_0:boot_flash_data_waitrequest
	wire  [14:0] mm_interconnect_0_boot_flash_data_address;                           // mm_interconnect_0:boot_flash_data_address -> boot_flash:avmm_data_addr
	wire         mm_interconnect_0_boot_flash_data_read;                              // mm_interconnect_0:boot_flash_data_read -> boot_flash:avmm_data_read
	wire         mm_interconnect_0_boot_flash_data_readdatavalid;                     // boot_flash:avmm_data_readdatavalid -> mm_interconnect_0:boot_flash_data_readdatavalid
	wire         mm_interconnect_0_boot_flash_data_write;                             // mm_interconnect_0:boot_flash_data_write -> boot_flash:avmm_data_write
	wire  [31:0] mm_interconnect_0_boot_flash_data_writedata;                         // mm_interconnect_0:boot_flash_data_writedata -> boot_flash:avmm_data_writedata
	wire   [1:0] mm_interconnect_0_boot_flash_data_burstcount;                        // mm_interconnect_0:boot_flash_data_burstcount -> boot_flash:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_e_debug_mem_slave_readdata;                  // nios2_e:debug_mem_slave_readdata -> mm_interconnect_0:nios2_e_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_waitrequest;               // nios2_e:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_e_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_debugaccess;               // mm_interconnect_0:nios2_e_debug_mem_slave_debugaccess -> nios2_e:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_e_debug_mem_slave_address;                   // mm_interconnect_0:nios2_e_debug_mem_slave_address -> nios2_e:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_read;                      // mm_interconnect_0:nios2_e_debug_mem_slave_read -> nios2_e:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_e_debug_mem_slave_byteenable;                // mm_interconnect_0:nios2_e_debug_mem_slave_byteenable -> nios2_e:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_write;                     // mm_interconnect_0:nios2_e_debug_mem_slave_write -> nios2_e:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_e_debug_mem_slave_writedata;                 // mm_interconnect_0:nios2_e_debug_mem_slave_writedata -> nios2_e:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                      // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                       // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                         // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                     // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                         // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_systimer_s1_chipselect;                            // mm_interconnect_0:systimer_s1_chipselect -> systimer:chipselect
	wire  [15:0] mm_interconnect_0_systimer_s1_readdata;                              // systimer:readdata -> mm_interconnect_0:systimer_s1_readdata
	wire   [2:0] mm_interconnect_0_systimer_s1_address;                               // mm_interconnect_0:systimer_s1_address -> systimer:address
	wire         mm_interconnect_0_systimer_s1_write;                                 // mm_interconnect_0:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_0_systimer_s1_writedata;                             // mm_interconnect_0:systimer_s1_writedata -> systimer:writedata
	wire         mm_interconnect_0_syskey_s1_chipselect;                              // mm_interconnect_0:syskey_s1_chipselect -> syskey:chipselect
	wire  [31:0] mm_interconnect_0_syskey_s1_readdata;                                // syskey:readdata -> mm_interconnect_0:syskey_s1_readdata
	wire   [1:0] mm_interconnect_0_syskey_s1_address;                                 // mm_interconnect_0:syskey_s1_address -> syskey:address
	wire         mm_interconnect_0_syskey_s1_write;                                   // mm_interconnect_0:syskey_s1_write -> syskey:write_n
	wire  [31:0] mm_interconnect_0_syskey_s1_writedata;                               // mm_interconnect_0:syskey_s1_writedata -> syskey:writedata
	wire         mm_interconnect_0_led7seg_s1_chipselect;                             // mm_interconnect_0:led7seg_s1_chipselect -> led7seg:chipselect
	wire  [31:0] mm_interconnect_0_led7seg_s1_readdata;                               // led7seg:readdata -> mm_interconnect_0:led7seg_s1_readdata
	wire   [1:0] mm_interconnect_0_led7seg_s1_address;                                // mm_interconnect_0:led7seg_s1_address -> led7seg:address
	wire         mm_interconnect_0_led7seg_s1_write;                                  // mm_interconnect_0:led7seg_s1_write -> led7seg:write_n
	wire  [31:0] mm_interconnect_0_led7seg_s1_writedata;                              // mm_interconnect_0:led7seg_s1_writedata -> led7seg:writedata
	wire         mm_interconnect_0_gpio_0_s1_chipselect;                              // mm_interconnect_0:gpio_0_s1_chipselect -> gpio_0:chipselect
	wire  [31:0] mm_interconnect_0_gpio_0_s1_readdata;                                // gpio_0:readdata -> mm_interconnect_0:gpio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_0_s1_address;                                 // mm_interconnect_0:gpio_0_s1_address -> gpio_0:address
	wire         mm_interconnect_0_gpio_0_s1_write;                                   // mm_interconnect_0:gpio_0_s1_write -> gpio_0:write_n
	wire  [31:0] mm_interconnect_0_gpio_0_s1_writedata;                               // mm_interconnect_0:gpio_0_s1_writedata -> gpio_0:writedata
	wire         mm_interconnect_0_gpio_1_s1_chipselect;                              // mm_interconnect_0:gpio_1_s1_chipselect -> gpio_1:chipselect
	wire  [31:0] mm_interconnect_0_gpio_1_s1_readdata;                                // gpio_1:readdata -> mm_interconnect_0:gpio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_1_s1_address;                                 // mm_interconnect_0:gpio_1_s1_address -> gpio_1:address
	wire         mm_interconnect_0_gpio_1_s1_write;                                   // mm_interconnect_0:gpio_1_s1_write -> gpio_1:write_n
	wire  [31:0] mm_interconnect_0_gpio_1_s1_writedata;                               // mm_interconnect_0:gpio_1_s1_writedata -> gpio_1:writedata
	wire         mm_interconnect_0_gpio_2_s1_chipselect;                              // mm_interconnect_0:gpio_2_s1_chipselect -> gpio_2:chipselect
	wire  [31:0] mm_interconnect_0_gpio_2_s1_readdata;                                // gpio_2:readdata -> mm_interconnect_0:gpio_2_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_2_s1_address;                                 // mm_interconnect_0:gpio_2_s1_address -> gpio_2:address
	wire         mm_interconnect_0_gpio_2_s1_write;                                   // mm_interconnect_0:gpio_2_s1_write -> gpio_2:write_n
	wire  [31:0] mm_interconnect_0_gpio_2_s1_writedata;                               // mm_interconnect_0:gpio_2_s1_writedata -> gpio_2:writedata
	wire         irq_mapper_receiver0_irq;                                            // systimer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                            // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_e_irq_irq;                                                     // irq_mapper:sender_irq -> nios2_e:irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [boot_flash:reset_n, gpio_0:reset_n, gpio_1:reset_n, gpio_2:reset_n, irq_mapper:reset, jtag_uart:rst_n, led7seg:reset_n, mm_interconnect_0:nios2_e_reset_reset_bridge_in_reset_reset, nios2_e:reset_n, onchip_memory2_0:reset, peridot_qspi_psram_0:csi_reset, rst_translator:in_reset, sysid:reset_n, syskey:reset_n, systimer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [nios2_e:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	altera_onchip_flash #(
		.INIT_FILENAME                       ("boot_onchip_flash.hex"),
		.INIT_FILENAME_SIM                   ("boot_onchip_flash.dat"),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M08SCE144C8G"),
		.DEVICE_ID                           ("08"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (23039),
		.SECTOR4_START_ADDR                  (0),
		.SECTOR4_END_ADDR                    (0),
		.SECTOR5_START_ADDR                  (0),
		.SECTOR5_END_ADDR                    (0),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (23039),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (23039),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (4),
		.SECTOR4_MAP                         (0),
		.SECTOR5_MAP                         (0),
		.ADDR_RANGE1_END_ADDR                (8191),
		.ADDR_RANGE2_END_ADDR                (23039),
		.ADDR_RANGE1_OFFSET                  (512),
		.ADDR_RANGE2_OFFSET                  (21504),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (15),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (2),
		.SECTOR_READ_PROTECTION_MODE         (24),
		.FLASH_SEQ_READ_DATA_COUNT           (2),
		.FLASH_ADDR_ALIGNMENT_BITS           (1),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (12),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (60),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (17500000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (15250),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) boot_flash (
		.clock                   (clk_clk),                                         //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                 // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_boot_flash_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_boot_flash_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_boot_flash_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_boot_flash_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_boot_flash_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_boot_flash_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_boot_flash_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_boot_flash_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_boot_flash_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_boot_flash_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_boot_flash_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_boot_flash_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_boot_flash_csr_readdata)        //       .readdata
	);

	nios2core_gpio_0 gpio_0 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_gpio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_0_s1_readdata),   //                    .readdata
		.bidir_port (gpio0_export)                            // external_connection.export
	);

	nios2core_gpio_0 gpio_1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_gpio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_1_s1_readdata),   //                    .readdata
		.bidir_port (gpio1_export)                            // external_connection.export
	);

	nios2core_gpio_0 gpio_2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_gpio_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_2_s1_readdata),   //                    .readdata
		.bidir_port (gpio2_export)                            // external_connection.export
	);

	nios2core_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	nios2core_led7seg led7seg (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led7seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led7seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led7seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led7seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led7seg_s1_readdata),   //                    .readdata
		.out_port   (led7seg_export)                           // external_connection.export
	);

	nios2core_nios2_e nios2_e (
		.clk                                 (clk_clk),                                               //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (nios2_e_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_e_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_e_data_master_read),                              //                          .read
		.d_readdata                          (nios2_e_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_e_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_e_data_master_write),                             //                          .write
		.d_writedata                         (nios2_e_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_e_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_e_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_e_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_e_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_e_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_e_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                      //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_e_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_e_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_e_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_e_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_e_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_e_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_e_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_e_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	nios2core_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	peridot_qspi_psram #(
		.CS_NEGATE_DELAY      (2),
		.CS_NEGATE_HOLD       (4),
		.SPI_READ_WAIT_CYCLE  (6),
		.QSPI_READ_WAIT_CYCLE (4),
		.READDATA_LATENCY     (4),
		.INITIAL_WAIT_CYCLE   (10),
		.DEVICE_FAMILY        ("MAX 10")
	) peridot_qspi_psram_0 (
		.avs_address       (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_address),       // avalon_slave_0.address
		.avs_read          (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_read),          //               .read
		.avs_readdata      (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_readdata),      //               .readdata
		.avs_readdatavalid (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_readdatavalid), //               .readdatavalid
		.avs_write         (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_write),         //               .write
		.avs_writedata     (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_writedata),     //               .writedata
		.avs_byteenable    (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_byteenable),    //               .byteenable
		.avs_waitrequest   (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_waitrequest),   //               .waitrequest
		.csi_reset         (rst_controller_reset_out_reset),                                      //     reset_sink.reset
		.csi_clock         (clk_clk),                                                             //     clock_sink.clk
		.qspi_sio          (qspi_sio),                                                            //    conduit_end.sio
		.qspi_sck          (qspi_sck),                                                            //               .sck
		.qspi_cs_n         (qspi_ce_n),                                                           //               .ce_n
		.outclock          (qspi_outclock)                                                        //               .outclock
	);

	nios2core_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	nios2core_syskey syskey (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_syskey_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_syskey_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_syskey_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_syskey_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_syskey_s1_readdata),   //                    .readdata
		.in_port    (syskey_in_port),                         // external_connection.export
		.out_port   (syskey_out_port)                         //                    .export
	);

	nios2core_systimer systimer (
		.clk        (clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_systimer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                  //   irq.irq
	);

	nios2core_mm_interconnect_0 mm_interconnect_0 (
		.clk_50m_clk_clk                                   (clk_clk),                                                             //                         clk_50m_clk.clk
		.nios2_e_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                      // nios2_e_reset_reset_bridge_in_reset.reset
		.nios2_e_data_master_address                       (nios2_e_data_master_address),                                         //                 nios2_e_data_master.address
		.nios2_e_data_master_waitrequest                   (nios2_e_data_master_waitrequest),                                     //                                    .waitrequest
		.nios2_e_data_master_byteenable                    (nios2_e_data_master_byteenable),                                      //                                    .byteenable
		.nios2_e_data_master_read                          (nios2_e_data_master_read),                                            //                                    .read
		.nios2_e_data_master_readdata                      (nios2_e_data_master_readdata),                                        //                                    .readdata
		.nios2_e_data_master_write                         (nios2_e_data_master_write),                                           //                                    .write
		.nios2_e_data_master_writedata                     (nios2_e_data_master_writedata),                                       //                                    .writedata
		.nios2_e_data_master_debugaccess                   (nios2_e_data_master_debugaccess),                                     //                                    .debugaccess
		.nios2_e_instruction_master_address                (nios2_e_instruction_master_address),                                  //          nios2_e_instruction_master.address
		.nios2_e_instruction_master_waitrequest            (nios2_e_instruction_master_waitrequest),                              //                                    .waitrequest
		.nios2_e_instruction_master_read                   (nios2_e_instruction_master_read),                                     //                                    .read
		.nios2_e_instruction_master_readdata               (nios2_e_instruction_master_readdata),                                 //                                    .readdata
		.boot_flash_csr_address                            (mm_interconnect_0_boot_flash_csr_address),                            //                      boot_flash_csr.address
		.boot_flash_csr_write                              (mm_interconnect_0_boot_flash_csr_write),                              //                                    .write
		.boot_flash_csr_read                               (mm_interconnect_0_boot_flash_csr_read),                               //                                    .read
		.boot_flash_csr_readdata                           (mm_interconnect_0_boot_flash_csr_readdata),                           //                                    .readdata
		.boot_flash_csr_writedata                          (mm_interconnect_0_boot_flash_csr_writedata),                          //                                    .writedata
		.boot_flash_data_address                           (mm_interconnect_0_boot_flash_data_address),                           //                     boot_flash_data.address
		.boot_flash_data_write                             (mm_interconnect_0_boot_flash_data_write),                             //                                    .write
		.boot_flash_data_read                              (mm_interconnect_0_boot_flash_data_read),                              //                                    .read
		.boot_flash_data_readdata                          (mm_interconnect_0_boot_flash_data_readdata),                          //                                    .readdata
		.boot_flash_data_writedata                         (mm_interconnect_0_boot_flash_data_writedata),                         //                                    .writedata
		.boot_flash_data_burstcount                        (mm_interconnect_0_boot_flash_data_burstcount),                        //                                    .burstcount
		.boot_flash_data_readdatavalid                     (mm_interconnect_0_boot_flash_data_readdatavalid),                     //                                    .readdatavalid
		.boot_flash_data_waitrequest                       (mm_interconnect_0_boot_flash_data_waitrequest),                       //                                    .waitrequest
		.gpio_0_s1_address                                 (mm_interconnect_0_gpio_0_s1_address),                                 //                           gpio_0_s1.address
		.gpio_0_s1_write                                   (mm_interconnect_0_gpio_0_s1_write),                                   //                                    .write
		.gpio_0_s1_readdata                                (mm_interconnect_0_gpio_0_s1_readdata),                                //                                    .readdata
		.gpio_0_s1_writedata                               (mm_interconnect_0_gpio_0_s1_writedata),                               //                                    .writedata
		.gpio_0_s1_chipselect                              (mm_interconnect_0_gpio_0_s1_chipselect),                              //                                    .chipselect
		.gpio_1_s1_address                                 (mm_interconnect_0_gpio_1_s1_address),                                 //                           gpio_1_s1.address
		.gpio_1_s1_write                                   (mm_interconnect_0_gpio_1_s1_write),                                   //                                    .write
		.gpio_1_s1_readdata                                (mm_interconnect_0_gpio_1_s1_readdata),                                //                                    .readdata
		.gpio_1_s1_writedata                               (mm_interconnect_0_gpio_1_s1_writedata),                               //                                    .writedata
		.gpio_1_s1_chipselect                              (mm_interconnect_0_gpio_1_s1_chipselect),                              //                                    .chipselect
		.gpio_2_s1_address                                 (mm_interconnect_0_gpio_2_s1_address),                                 //                           gpio_2_s1.address
		.gpio_2_s1_write                                   (mm_interconnect_0_gpio_2_s1_write),                                   //                                    .write
		.gpio_2_s1_readdata                                (mm_interconnect_0_gpio_2_s1_readdata),                                //                                    .readdata
		.gpio_2_s1_writedata                               (mm_interconnect_0_gpio_2_s1_writedata),                               //                                    .writedata
		.gpio_2_s1_chipselect                              (mm_interconnect_0_gpio_2_s1_chipselect),                              //                                    .chipselect
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),               //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                 //                                    .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                  //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),              //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),             //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),           //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),            //                                    .chipselect
		.led7seg_s1_address                                (mm_interconnect_0_led7seg_s1_address),                                //                          led7seg_s1.address
		.led7seg_s1_write                                  (mm_interconnect_0_led7seg_s1_write),                                  //                                    .write
		.led7seg_s1_readdata                               (mm_interconnect_0_led7seg_s1_readdata),                               //                                    .readdata
		.led7seg_s1_writedata                              (mm_interconnect_0_led7seg_s1_writedata),                              //                                    .writedata
		.led7seg_s1_chipselect                             (mm_interconnect_0_led7seg_s1_chipselect),                             //                                    .chipselect
		.nios2_e_debug_mem_slave_address                   (mm_interconnect_0_nios2_e_debug_mem_slave_address),                   //             nios2_e_debug_mem_slave.address
		.nios2_e_debug_mem_slave_write                     (mm_interconnect_0_nios2_e_debug_mem_slave_write),                     //                                    .write
		.nios2_e_debug_mem_slave_read                      (mm_interconnect_0_nios2_e_debug_mem_slave_read),                      //                                    .read
		.nios2_e_debug_mem_slave_readdata                  (mm_interconnect_0_nios2_e_debug_mem_slave_readdata),                  //                                    .readdata
		.nios2_e_debug_mem_slave_writedata                 (mm_interconnect_0_nios2_e_debug_mem_slave_writedata),                 //                                    .writedata
		.nios2_e_debug_mem_slave_byteenable                (mm_interconnect_0_nios2_e_debug_mem_slave_byteenable),                //                                    .byteenable
		.nios2_e_debug_mem_slave_waitrequest               (mm_interconnect_0_nios2_e_debug_mem_slave_waitrequest),               //                                    .waitrequest
		.nios2_e_debug_mem_slave_debugaccess               (mm_interconnect_0_nios2_e_debug_mem_slave_debugaccess),               //                                    .debugaccess
		.onchip_memory2_0_s1_address                       (mm_interconnect_0_onchip_memory2_0_s1_address),                       //                 onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                         (mm_interconnect_0_onchip_memory2_0_s1_write),                         //                                    .write
		.onchip_memory2_0_s1_readdata                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                      //                                    .readdata
		.onchip_memory2_0_s1_writedata                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                     //                                    .writedata
		.onchip_memory2_0_s1_byteenable                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                    //                                    .byteenable
		.onchip_memory2_0_s1_chipselect                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                    //                                    .chipselect
		.onchip_memory2_0_s1_clken                         (mm_interconnect_0_onchip_memory2_0_s1_clken),                         //                                    .clken
		.peridot_qspi_psram_0_avalon_slave_0_address       (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_address),       // peridot_qspi_psram_0_avalon_slave_0.address
		.peridot_qspi_psram_0_avalon_slave_0_write         (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_write),         //                                    .write
		.peridot_qspi_psram_0_avalon_slave_0_read          (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_read),          //                                    .read
		.peridot_qspi_psram_0_avalon_slave_0_readdata      (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_readdata),      //                                    .readdata
		.peridot_qspi_psram_0_avalon_slave_0_writedata     (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_writedata),     //                                    .writedata
		.peridot_qspi_psram_0_avalon_slave_0_byteenable    (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_byteenable),    //                                    .byteenable
		.peridot_qspi_psram_0_avalon_slave_0_readdatavalid (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_readdatavalid), //                                    .readdatavalid
		.peridot_qspi_psram_0_avalon_slave_0_waitrequest   (mm_interconnect_0_peridot_qspi_psram_0_avalon_slave_0_waitrequest),   //                                    .waitrequest
		.sysid_control_slave_address                       (mm_interconnect_0_sysid_control_slave_address),                       //                 sysid_control_slave.address
		.sysid_control_slave_readdata                      (mm_interconnect_0_sysid_control_slave_readdata),                      //                                    .readdata
		.syskey_s1_address                                 (mm_interconnect_0_syskey_s1_address),                                 //                           syskey_s1.address
		.syskey_s1_write                                   (mm_interconnect_0_syskey_s1_write),                                   //                                    .write
		.syskey_s1_readdata                                (mm_interconnect_0_syskey_s1_readdata),                                //                                    .readdata
		.syskey_s1_writedata                               (mm_interconnect_0_syskey_s1_writedata),                               //                                    .writedata
		.syskey_s1_chipselect                              (mm_interconnect_0_syskey_s1_chipselect),                              //                                    .chipselect
		.systimer_s1_address                               (mm_interconnect_0_systimer_s1_address),                               //                         systimer_s1.address
		.systimer_s1_write                                 (mm_interconnect_0_systimer_s1_write),                                 //                                    .write
		.systimer_s1_readdata                              (mm_interconnect_0_systimer_s1_readdata),                              //                                    .readdata
		.systimer_s1_writedata                             (mm_interconnect_0_systimer_s1_writedata),                             //                                    .writedata
		.systimer_s1_chipselect                            (mm_interconnect_0_systimer_s1_chipselect)                             //                                    .chipselect
	);

	nios2core_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_e_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
